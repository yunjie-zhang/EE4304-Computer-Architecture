module Decoder(in, out);
    parameter WORD = 32;

    input [4:0] in;

    output reg [WORD - 1:0] out;


    always @* begin
        case(in)
            5'b00000: out <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
            5'b00001: out <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
            5'b00010: out <= 32'b0000_0000_0000_0000_0000_0000_0000_0100;
            5'b00011: out <= 32'b0000_0000_0000_0000_0000_0000_0000_1000;
            5'b00100: out <= 32'b0000_0000_0000_0000_0000_0000_0001_0000;
            5'b00101: out <= 32'b0000_0000_0000_0000_0000_0000_0010_0000;
            5'b00110: out <= 32'b0000_0000_0000_0000_0000_0000_0100_0000;
            5'b00111: out <= 32'b0000_0000_0000_0000_0000_0000_1000_0000;
            5'b01000: out <= 32'b0000_0000_0000_0000_0000_0001_0000_0000;
            5'b01001: out <= 32'b0000_0000_0000_0000_0000_0010_0000_0000;
            5'b01010: out <= 32'b0000_0000_0000_0000_0000_0100_0000_0000;
            5'b01011: out <= 32'b0000_0000_0000_0000_0000_1000_0000_0000;
            5'b01100: out <= 32'b0000_0000_0000_0000_0001_0000_0000_0000;
            5'b01101: out <= 32'b0000_0000_0000_0000_0010_0000_0000_0000;
            5'b01110: out <= 32'b0000_0000_0000_0000_0100_0000_0000_0000;
            5'b01111: out <= 32'b0000_0000_0000_0000_1000_0000_0000_0000;
            5'b10000: out <= 32'b0000_0000_0000_0001_0000_0000_0000_0000;
            5'b10001: out <= 32'b0000_0000_0000_0010_0000_0000_0000_0000;
            5'b10010: out <= 32'b0000_0000_0000_0100_0000_0000_0000_0000;
            5'b10011: out <= 32'b0000_0000_0000_1000_0000_0000_0000_0000;
            5'b10100: out <= 32'b0000_0000_0001_0000_0000_0000_0000_0000;
            5'b10101: out <= 32'b0000_0000_0010_0000_0000_0000_0000_0000;
            5'b10110: out <= 32'b0000_0000_0100_0000_0000_0000_0000_0000;
            5'b10111: out <= 32'b0000_0000_1000_0000_0000_0000_0000_0000;
            5'b11000: out <= 32'b0000_0001_0000_0000_0000_0000_0000_0000;
            5'b11001: out <= 32'b0000_0010_0000_0000_0000_0000_0000_0000;
            5'b11010: out <= 32'b0000_0100_0000_0000_0000_0000_0000_0000;
            5'b11011: out <= 32'b0000_1000_0000_0000_0000_0000_0000_0000;
            5'b11100: out <= 32'b0001_0000_0000_0000_0000_0000_0000_0000;
            5'b11101: out <= 32'b0010_0000_0000_0000_0000_0000_0000_0000;
            5'b11110: out <= 32'b0100_0000_0000_0000_0000_0000_0000_0000;
            5'b11111: out <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
        endcase
    end

endmodule
